* Created by KLayout

* cell bgr_simple
.SUBCKT bgr_simple
* net 1 Vout
* net 2 Vin
* net 26 Gnd
* device instance $4 r0 *1 -75.5,-147.5 RES
R$4 10 26 28800
* device instance $16 r0 *1 -27.5,-147.5 RES
R$16 25 10 4000
* device instance $75 r0 *1 86.6,-59.5 RES
R$75 13 3 28000
* device instance $97 r0 *1 44.4,-25.9 RES
R$97 3 1 1000
* device instance $98 r0 *1 59.5,-80 HRES
R$98 7 2 1050000
* device instance $102 r0 *1 24.3,-65.2 NMOS
M$102 3 7 7 26 NMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $104 r0 *1 6.3,-65.2 NMOS
M$104 8 7 6 26 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $105 r0 *1 15.3,-65.2 NMOS
M$105 11 7 9 26 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $106 r0 *1 15.3,-28 PMOS
M$106 2 6 9 2 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $107 r0 *1 6.3,-28 PMOS
M$107 2 6 6 2 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $108 r0 *1 24.3,-28 PMOS
M$108 2 9 7 2 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $110 r180 *1 52.2,-173.5 PMOS
M$110 13 13 13 26 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $112 r180 *1 36.7,-96.5 PMOS
M$112 11 11 11 25 PMOS L=1U W=160U AS=320P AD=320P PS=352U PD=352U
* device instance $120 r180 *1 23.2,-134 PMOS
M$120 8 8 8 10 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS bgr_simple
