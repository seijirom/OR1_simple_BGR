* Created by KLayout

* cell bgr_simple
.SUBCKT bgr_simple
* net 1 Vin
* net 4 R2
* net 5 R1
* net 9 Rex
* net 11 R3
* net 13 D
* net 26 Gnd
* device instance $1 r270 *1 27,-47.5 D
D$1 26 6 D A=4P P=8U
* device instance $2 r90 *1 2.5,-48.5 D
D$2 26 7 D A=4P P=8U
* device instance $3 m45 *1 12.5,-48.5 D
D$3 26 10 D A=4P P=8U
* device instance $4 r180 *1 52.5,-21.5 RES
R$4 12 3 1000 RES
* device instance $11 r180 *1 47.5,-80 HRES
R$11 6 9 1050000 HRES
* device instance $15 m90 *1 90.5,-59.5 RES
R$15 13 3 28000 RES
* device instance $40 m90 *1 -20,-147.5 RES
R$40 25 8 4000 RES
* device instance $81 m90 *1 -36,-147.5 RES
R$81 8 26 25600 RES
* device instance $100 r0 *1 6,-65.5 NMOS
M$100 2 6 7 26 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $101 r0 *1 24,-65.5 NMOS
M$101 3 6 6 26 NMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $103 r0 *1 15,-65.5 NMOS
M$103 20 6 10 26 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $104 r0 *1 15.5,-27.5 PMOS
M$104 1 7 10 1 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $105 r0 *1 24.5,-27.5 PMOS
M$105 1 10 6 1 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $106 r0 *1 6.5,-27.5 PMOS
M$106 1 7 7 1 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $108 r180 *1 52,-174 PMOS
M$108 13 13 13 26 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $110 r180 *1 36.5,-97 PMOS
M$110 20 20 20 25 PMOS L=1U W=160U AS=320P AD=320P PS=352U PD=352U
* device instance $118 r180 *1 23,-134.5 PMOS
M$118 2 2 2 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS bgr_simple
