* Created by KLayout

* cell bgr_simple
* pin Vin
* pin R2
* pin R1
* pin Rex
* pin R3
* pin Vout
* pin D
* pin Gnd
.SUBCKT bgr_simple 2 4 5 8 11 12 13 26
* net 2 Vin
* net 4 R2
* net 5 R1
* net 8 Rex
* net 11 R3
* net 12 Vout
* net 13 D
* net 26 Gnd
* device instance $1 m0 *1 58.5,-72.5 HRES
R$1 8 6 1050000 HRES
* device instance $6 r270 *1 27,-47.5 D
D$6 26 6 D A=4P P=8U
* device instance $7 r90 *1 2.5,-48.5 D
D$7 26 7 D A=4P P=8U
* device instance $8 m45 *1 12.5,-48.5 D
D$8 26 10 D A=4P P=8U
* device instance $9 r180 *1 52.5,-21.5 RES
R$9 12 3 1000 RES
* device instance $16 m90 *1 90.5,-59.5 RES
R$16 5 3 2000 RES
* device instance $26 m90 *1 150.5,-59.5 RES
R$26 11 4 4000 RES
* device instance $31 m90 *1 110.5,-59.5 RES
R$31 5 4 2000 RES
* device instance $41 m90 *1 -20,-147.5 RES
R$41 25 9 4000 RES
* device instance $82 m90 *1 -36,-147.5 RES
R$82 9 26 25600 RES
* device instance $97 m90 *1 94.5,-147.5 RES
R$97 13 11 20000 RES
* device instance $101 r0 *1 6,-65.5 NMOS
M$101 1 6 7 26 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $102 r0 *1 33,-65.5 NMOS
M$102 3 6 6 26 NMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $104 r0 *1 15,-65.5 NMOS
M$104 20 6 10 26 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $105 r0 *1 15.5,-27.5 PMOS
M$105 2 7 10 2 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $106 r0 *1 24.5,-27.5 PMOS
M$106 2 10 6 2 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $107 r0 *1 6.5,-27.5 PMOS
M$107 2 7 7 2 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $109 r180 *1 52,-174 PMOS
M$109 13 13 13 26 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $111 r180 *1 36.5,-97 PMOS
M$111 20 20 20 25 PMOS L=1U W=160U AS=320P AD=320P PS=352U PD=352U
* device instance $119 r180 *1 22.5,-134.5 PMOS
M$119 1 1 1 9 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS bgr_simple
