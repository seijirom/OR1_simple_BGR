* Z:\HOME\SEIJIROM\WORK\2021_9\OR1_SIMPLE_BGR\BGR_SIMPLE_TB.ASC
*V1 N001 0 5
R1 N002 0 1MEG
XX1 N001 N002 N001 N003 N004 N005 N006 BGR_SIMPLE

* BLOCK SYMBOL DEFINITIONS
.SUBCKT BGR_SIMPLE VIN VOUT REX D R1 R2 R3
M1 N003 N002 VIN VIN PMOS L=1U W=40U
M2 N002 N001 VIN VIN PMOS L=1U W=20U
M3 N001 N001 VIN VIN PMOS L=1U W=20U
M4 N003 N003 N004 0 NMOS L=1U W=40U
M5 N002 N003 N006 0 NMOS L=1U W=20U
M6 N001 N003 N005 0 NMOS L=1U W=20U
R1 REX N003 1.005MEG
R2 N008 N012 4K
R5 VOUT N004 1K
M7 N005 N005 N005 N012 PMOS L=1U W=20U
M8 N006 N006 N006 N008 PMOS L=1U W=160U
M9 D D D 0 PMOS L=1U W=40U
D1 0 N001 D
D2 0 N002 D
D4 0 N003 D
R3 N007 N010 4K
R4 N010 N013 4K
R6 N013 N012 1.6K
R7 N007 N011 4K
R8 N011 N014 4K
R9 N014 N016 4K
R10 N016 0 4K
R11 N018 N017 4K
R12 N017 N015 4K
R13 N015 N009 4K
R14 N018 R3 4K
R15 R3 R2 4K
R16 R2 R1 4K
R17 R1 N004 4K
R18 D N009 4K
R20 R1 N004 4K
R21 R2 R1 4K
.ENDS BGR_SIMPLE

.MODEL D D
.LIB C:\USERS\SEIJIROM\MY DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.DIO
.MODEL NMOS NMOS
.MODEL PMOS PMOS
.LIB C:\USERS\SEIJIROM\MY DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.MOS
* .STEP PARAM R LIST   29.6K 29.7K 29.8K 29.9K 30K 30.1K
.DC TEMP _40 120 1
.PARAM R=29.8K
*.INCLUDE "./MODELS/OR1_MOS"
* .AC DEC 1 1 10
.BACKANNO
.GLOBAL 0
.END
