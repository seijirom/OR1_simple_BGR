* Created by KLayout

* cell bgr_simple
.SUBCKT bgr_simple
* net 8 SUBSTRATE
* device instance $1 r0 *1 -87.5,-147.5 RES
R$1 2 2 40
* device instance $16 r0 *1 -27.5,-147.5 RES
R$16 6 6 38.0952380952
* device instance $21 r0 *1 166.5,-147.5 RES
R$21 1 1 16
* device instance $46 r0 *1 59.5,-80 RES
R$46 9 9 187.5
* device instance $96 r0 *1 59.5,-80 HRES
R$96 9 9 65625
* device instance $100 r0 *1 6.3,-65.2 NMOS
M$100 8 5 3 8 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $101 r0 *1 33.3,-65.2 NMOS
M$101 8 5 4 8 NMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $103 r0 *1 15.3,-65.2 NMOS
M$103 8 5 5 8 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $104 r0 *1 6.3,-28 PMOS
M$104 7 3 3 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $105 r0 *1 15.3,-28 PMOS
M$105 7 3 5 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $106 r0 *1 33.3,-28 PMOS
M$106 7 5 4 7 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $108 r180 *1 52.2,-173.5 PMOS
M$108 1 1 1 2 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $110 r180 *1 36.7,-96.5 PMOS
M$110 8 8 8 6 PMOS L=1U W=180U AS=360P AD=360P PS=396U PD=396U
.ENDS bgr_simple
