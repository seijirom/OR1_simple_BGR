* Created by KLayout

* cell bgr_simple
.SUBCKT bgr_simple
* net 1 Vout
* net 2 Vin
* net 5 R2
* net 6 R1
* net 11 D
* net 12 R3
* net 26 Gnd
* device instance $19 r0 *1 -15.5,-147.5 RES
R$19 9 25 4000
* device instance $61 r0 *1 -27.5,-59.5 RES
R$61 9 26 28800
* device instance $79 r0 *1 86.5,-59.5 RES
R$79 11 4 28000
* device instance $93 r0 *1 60.5,-21.5 RES
R$93 4 1 1000
* device instance $97 r0 *1 59.5,-80 HRES
R$97 7 2 1050000
* device instance $101 r270 *1 27,-47.5 D
D$101 26 106 D A=1P P=4U
* device instance $102 r90 *1 2.5,-48.5 D
D$102 26 107 D A=1P P=4U
* device instance $103 m45 *1 12.5,-48.5 D
D$103 26 108 D A=1P P=4U
* device instance $104 r0 *1 6,-65.5 NMOS
M$104 3 7 8 26 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $105 r0 *1 24,-65.5 NMOS
M$105 4 7 7 26 NMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $107 r0 *1 15,-65.5 NMOS
M$107 13 7 10 26 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $108 r0 *1 15.5,-27.5 PMOS
M$108 2 8 10 2 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $109 r0 *1 6.5,-27.5 PMOS
M$109 2 8 8 2 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $110 r0 *1 24.5,-27.5 PMOS
M$110 2 10 7 2 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $112 r180 *1 52,-174 PMOS
M$112 11 11 11 26 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $114 r180 *1 36.5,-97 PMOS
M$114 13 13 13 25 PMOS L=1U W=160U AS=320P AD=320P PS=352U PD=352U
* device instance $122 r180 *1 23,-134.5 PMOS
M$122 3 3 3 9 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS bgr_simple
