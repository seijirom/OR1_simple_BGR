* Created by KLayout

* cell bgr_simple
.SUBCKT bgr_simple
* net 1 Vout
* net 2 Vin
* net 5 R2
* net 6 R1
* net 11 D
* net 12 R3
* net 25 Gnd
* cell instance $1 r180 *1 65.5,-10
X$1 4 1 R_poly$2
* cell instance $2 r180 *1 60.5,-41
X$2 2 7 HR_poly
* cell instance $3 r0 *1 12,-43
X$3 2 8 10 2 pch1x20
* cell instance $4 r0 *1 21,-43
X$4 2 10 7 2 pch1x20
* cell instance $5 r0 *1 3,-43
X$5 2 8 8 2 pch1x20
* cell instance $6 r0 *1 30,-43
X$6 2 10 7 2 pch1x20
* cell instance $7 r0 *1 3,-78
X$7 25 7 8 3 nch1x20
* cell instance $8 r180 *1 39.5,-151.5
X$8 19 24 9 3 diodeblock
* cell instance $9 m90 *1 107.5,-101
X$9 6 4 R_poly$5
* cell instance $10 r0 *1 69.5,-101
X$10 6 4 R_poly$5
* cell instance $11 r0 *1 21,-78
X$11 25 7 7 4 nch1x20
* cell instance $12 r0 *1 30,-78
X$12 25 7 7 4 nch1x20
* cell instance $13 m90 *1 127.5,-101
X$13 6 5 R_poly$5
* cell instance $14 m90 *1 167.5,-101
X$14 12 5 R_poly$5
* cell instance $15 r0 *1 129.5,-101
X$15 6 5 R_poly$5
* cell instance $16 r0 *1 12,-78
X$16 25 7 10 19 nch1x20
* cell instance $17 r270 *1 3,-43
X$17 25 protection
* cell instance $18 r90 *1 26.5,-53
X$18 25 protection
* cell instance $19 r180 *1 -15,-18
X$19 9 14 R_poly
* cell instance $20 m90 *1 -3,-189
X$20 24 9 R_poly$5
* cell instance $21 m45 *1 -11.5,-53
X$21 25 protection
* cell instance $22 r0 *1 69.5,-189
X$22 11 20 R_poly$5
* cell instance $23 r180 *1 57.5,-123
X$23 11 25 pchdiode
* cell instance $24 r180 *1 57.5,-157.5
X$24 11 25 pchdiode
* cell instance $25 r0 *1 149.5,-189
X$25 23 12 R_poly$5
* cell instance $26 m0 *1 -61,-18
X$26 13 15 R_poly$5
* cell instance $27 r180 *1 -63,-18
X$27 13 16 R_poly$5
* cell instance $28 r180 *1 -23,-18
X$28 14 15 R_poly$5
* cell instance $29 m90 *1 -63,-189
X$29 17 16 R_poly$5
* cell instance $30 r0 *1 -61,-189
X$30 17 18 R_poly$5
* cell instance $31 m90 *1 -23,-189
X$31 25 18 R_poly$5
* cell instance $32 m90 *1 107.5,-189
X$32 21 20 R_poly$5
* cell instance $33 r0 *1 109.5,-189
X$33 21 22 R_poly$5
* cell instance $34 m90 *1 147.5,-189
X$34 23 22 R_poly$5
.ENDS bgr_simple

* cell protection
* pin 
.SUBCKT protection 2
* device instance $1 r0 *1 4.5,24 D
D$1 2 1 D A=1P P=4U
.ENDS protection

* cell R_poly$2
* pin 
* pin 
.SUBCKT R_poly$2 5 6
* device instance $1 r0 *1 13,11.5 RES
R$1 4 3 200 RES
* device instance $2 r0 *1 17,11.5 RES
R$2 4 6 200 RES
* device instance $3 r0 *1 9,11.5 RES
R$3 2 3 200 RES
* device instance $4 r0 *1 5,11.5 RES
R$4 2 1 200 RES
* device instance $5 r0 *1 1,11.5 RES
R$5 5 1 200 RES
.ENDS R_poly$2

* cell R_poly
* pin 
* pin 
.SUBCKT R_poly 2 3
* device instance $1 r0 *1 5,41.5 RES
R$1 3 1 800 RES
* device instance $2 r0 *1 1,41.5 RES
R$2 2 1 800 RES
.ENDS R_poly

* cell HR_poly
* pin 
* pin 
.SUBCKT HR_poly 4 5
* device instance $1 r0 *1 13,39 HRES
R$1 5 3 262500 HRES
* device instance $2 r0 *1 9,39 HRES
R$2 2 3 262500 HRES
* device instance $3 r0 *1 5,39 HRES
R$3 2 1 262500 HRES
* device instance $4 r0 *1 1,39 HRES
R$4 4 1 262500 HRES
.ENDS HR_poly

* cell R_poly$5
* pin 
* pin 
.SUBCKT R_poly$5 5 6
* device instance $1 r0 *1 17,41.5 RES
R$1 4 6 800 RES
* device instance $2 r0 *1 13,41.5 RES
R$2 4 3 800 RES
* device instance $3 r0 *1 9,41.5 RES
R$3 2 3 800 RES
* device instance $4 r0 *1 5,41.5 RES
R$4 2 1 800 RES
* device instance $5 r0 *1 1,41.5 RES
R$5 5 1 800 RES
.ENDS R_poly$5

* cell diodeblock
* pin 
* pin 
* pin 
* pin 
.SUBCKT diodeblock 1 2 3 4
* cell instance $1 r0 *1 -2.5,-71
X$1 1 2 pchdiode
* cell instance $2 r0 *1 25.5,-71
X$2 1 2 pchdiode
* cell instance $3 r0 *1 11,-71
X$3 1 2 pchdiode
* cell instance $4 r0 *1 25.5,-33.5
X$4 1 2 pchdiode
* cell instance $5 r0 *1 -2.5,-33.5
X$5 1 2 pchdiode
* cell instance $6 r0 *1 25.5,4
X$6 1 2 pchdiode
* cell instance $7 r0 *1 11,4
X$7 1 2 pchdiode
* cell instance $8 r0 *1 -2.5,4
X$8 1 2 pchdiode
* cell instance $9 r0 *1 11,-33.5
X$9 4 3 pchdiode
.ENDS diodeblock

* cell nch1x20
* pin SUBSTRATE
* pin 
* pin 
* pin 
.SUBCKT nch1x20 1 2 3 4
* net 1 SUBSTRATE
* cell instance $1 r0 *1 0.5,-0.5
X$1 4 3 2 1 Nch
.ENDS nch1x20

* cell Nch
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 2.5,13 NMOS
M$1 1 3 2 4 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS Nch

* cell pchdiode
* pin 
* pin 
.SUBCKT pchdiode 1 2
* cell instance $1 r0 *1 2,1
X$1 2 1 1 1 pch1x20
.ENDS pchdiode

* cell pch1x20
* pin 
* pin 
* pin 
* pin 
.SUBCKT pch1x20 1 2 3 4
* cell instance $1 r0 *1 1,2.5
X$1 4 3 2 1 Pch
.ENDS pch1x20

* cell Pch
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch 1 2 3 4
* device instance $1 r0 *1 2.5,13 PMOS
M$1 1 3 2 4 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS Pch
