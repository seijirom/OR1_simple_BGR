* C:\USERS\SEIJIROM\DROPBOX\MAKELSI\2020T^9G\BGR\BGR_SIMPLE_TB.ASC
*V1 N001 0 5
*R1 N002 0 1MEG
XX1 N001 N002 BGR_SIMPLE

* BLOCK SYMBOL DEFINITIONS
.SUBCKT BGR_SIMPLE VIN VOUT
M1 N003 N002 VIN VIN PCH L=1U W=40.0U M=1
M2 N002 N001 VIN VIN PCH L=1U W=20U
M3 N001 N001 VIN VIN PCH L=1U W=20U
M4 N003 N003 N004 0 NCH L=1U W=40.0U M=1
M5 N002 N003 N006 0 NCH L=1U W=20U
M6 N001 N003 N005 0 NCH L=1U W=20U
R1 VIN N003 1.005MEG
R2 N008 N013 4K
R5 VOUT N004 1K

M7 N005 N005 N005 N013 PCH L=1U W=20U
M8 N006 N006 N006 N008 PCH L=1U W=160U
M9 N018 N018 N018 0 PCH L=1U W=40U
D1 0 N001 D
D2 0 N002 D
D3 0 N004 D
D4 0 N003 D
R3 N007 N010 4K
R4 N010 N014 4K
R6 N014 N022 4K
R7 N007 N011 4K
R8 N011 N015 4K
R9 N015 N021 4K
R10 N021 0 4K
R11 N023 N019 4K
R12 N019 N016 4K
R13 N016 N009 4K
R14 N023 N020 4K
R15 N020 N017 4K
R16 N017 N012 2K
R17 N012 N004 2K
R18 N018 N009 4K
R19 N022 N013 800
.ENDS BGR_SIMPLE

.MODEL D D
.LIB C:\USERS\SEIJIROM\DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.DIO
.MODEL NMOS NMOS
.MODEL PMOS PMOS
.LIB C:\USERS\SEIJIROM\DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.MOS
* .STEP PARAM R LIST   29.6K 29.7K 29.8K 29.9K 30K 30.1K
.DC TEMP _40 120 1
.PARAM R=29.8K
*.INCLUDE "./MODELS/OR1_MOS"
.BACKANNO
.END
